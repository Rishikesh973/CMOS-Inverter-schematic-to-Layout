magic
tech sky130A
timestamp 1695408433
<< nwell >>
rect 450 350 750 815
<< nmos >>
rect 595 35 610 165
<< pmos >>
rect 595 395 610 605
<< ndiff >>
rect 540 155 595 165
rect 540 45 550 155
rect 580 45 595 155
rect 540 35 595 45
rect 610 155 665 165
rect 610 45 625 155
rect 655 45 665 155
rect 610 35 665 45
<< pdiff >>
rect 550 595 595 605
rect 550 405 560 595
rect 585 405 595 595
rect 550 395 595 405
rect 610 595 655 605
rect 610 405 625 595
rect 650 405 655 595
rect 610 395 655 405
<< ndiffc >>
rect 550 45 580 155
rect 625 45 655 155
<< pdiffc >>
rect 560 405 585 595
rect 625 405 650 595
<< psubdiff >>
rect 545 -10 660 5
rect 545 -35 560 -10
rect 635 -35 660 -10
rect 545 -50 660 -35
<< nsubdiff >>
rect 545 775 660 795
rect 545 750 560 775
rect 645 750 660 775
rect 545 735 660 750
<< psubdiffcont >>
rect 560 -35 635 -10
<< nsubdiffcont >>
rect 560 750 645 775
<< poly >>
rect 595 605 610 700
rect 595 355 610 395
rect 545 345 610 355
rect 545 325 555 345
rect 575 325 610 345
rect 545 315 610 325
rect 670 345 705 355
rect 670 325 680 345
rect 700 325 705 345
rect 670 315 705 325
rect 595 165 610 315
rect 595 20 610 35
<< polycont >>
rect 555 325 575 345
rect 680 325 700 345
<< locali >>
rect 545 775 660 795
rect 545 750 560 775
rect 645 750 660 775
rect 545 735 660 750
rect 550 595 595 735
rect 550 405 560 595
rect 585 575 595 595
rect 615 595 655 605
rect 585 405 590 575
rect 550 395 590 405
rect 615 405 625 595
rect 650 405 655 595
rect 615 395 655 405
rect 625 355 650 395
rect 545 345 580 355
rect 545 325 555 345
rect 575 325 580 345
rect 545 315 580 325
rect 625 345 705 355
rect 625 325 680 345
rect 700 325 705 345
rect 625 315 705 325
rect 625 165 650 315
rect 540 155 590 165
rect 540 45 550 155
rect 580 45 590 155
rect 540 35 590 45
rect 615 155 665 165
rect 615 45 625 155
rect 655 45 665 155
rect 615 35 665 45
rect 540 5 580 35
rect 540 -10 660 5
rect 540 -35 560 -10
rect 635 -35 660 -10
rect 540 -45 660 -35
rect 545 -50 660 -45
<< viali >>
rect 590 750 615 775
rect 585 -35 610 -10
<< metal1 >>
rect 270 775 995 800
rect 270 750 590 775
rect 615 750 995 775
rect 270 725 995 750
rect 450 315 580 355
rect 625 315 855 355
rect 265 -10 990 15
rect 265 -35 585 -10
rect 610 -35 990 -10
rect 265 -60 990 -35
<< labels >>
rlabel metal1 820 755 820 755 1 vdd
rlabel metal1 800 -20 800 -20 1 vss
rlabel metal1 770 330 780 340 1 out
rlabel metal1 490 325 500 335 1 in
<< end >>
