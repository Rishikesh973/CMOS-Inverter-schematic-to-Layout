* SPICE3 file created from inv_layout.ext - technology: sky130A

X0 a_1220_70# a_1090_630# vss vss sky130_fd_pr__nfet_01v8 ad=0.715 pd=3.7 as=0.715 ps=3.7 w=1.3 l=0.15
X1 a_1220_70# a_1090_630# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.945 pd=5.1 as=0.945 ps=5.1 w=2.1 l=0.15
C0 vdd vss 2.41f **FLOATING
