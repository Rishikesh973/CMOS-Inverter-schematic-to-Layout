** sch_path: /home/rishikesh/Desktop/cmos_inv/inverter_TB.sch
**.subckt inverter_TB
Vin vin GND PULSE(0 1.8 0 0.1n 0.1n 10n 20n 10)
.save i(vin)
vdd vdd GND 1.8
.save i(vdd)
x1 vdd vin vout GND inverter_vtc
C1 vout GND 0.5p m=1
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.dc vin 0 2 1m
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  inverter_vtc.sym # of pins=4
** sym_path: /home/rishikesh/Desktop/cmos_inv/inverter_vtc.sym
** sch_path: /home/rishikesh/Desktop/cmos_inv/inverter_vtc.sch
.subckt inverter_vtc vdd vin vout gnd
*.ipin vin
*.ipin gnd
*.opin vout
*.ipin vdd
XM1 vout vin gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
